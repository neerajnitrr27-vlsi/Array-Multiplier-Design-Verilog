`timescale 1ns / 1ps

// ---------------- Half Adder ----------------
module ha(
    input a, b,
    output sum, carry
);
    assign sum = a ^ b;
    assign carry = a & b;
endmodule

// ---------------- Full Adder ----------------
module fa (
    input a, b, cin,
    output sum, carry
);
    assign sum = a ^ b ^ cin;
    assign carry = (a & b) | (b & cin) | (a & cin);
endmodule

// ---------------- 32x32  Multiplier ----------------
module multi_32bit (
    input [31:0] A, B,
    output [63:0] m
);
    wire [1023:0] p;
    wire [2046:0] s, c;

    genvar i, j;

    // Generate Partial Products
    generate
        for(j = 0; j < 32; j = j + 1) begin: row
            for(i = 0; i < 32; i = i + 1) begin: col
                assign p[i + j*32] = A[i] & B[j];
            end
        end
    endgenerate



ha ha0(p[1], p[32], s[0], c[0]);

fa fa0(p[2], p[33], c[0], s[1], c[1]);
ha ha1(p[64], s[1], s[2], c[2]);

fa fa1(p[3], p[34], c[1], s[3], c[3]);
fa fa2(p[65], s[3], c[2], s[4], c[4]);
ha ha2(p[96], s[4], s[5], c[5]);

fa fa3(p[4], p[35], c[3], s[6], c[6]);
fa fa4(p[66], s[6], c[4], s[7], c[7]);
fa fa5(p[97], s[7], c[5], s[8], c[8]);
ha ha3(p[128], s[8], s[9], c[9]);

fa fa6(p[5], p[36], c[6], s[10], c[10]);
fa fa7(p[67], s[10], c[7], s[11], c[11]);
fa fa8(p[98], s[11], c[8], s[12], c[12]);
fa fa9(p[129], s[12], c[9], s[13], c[13]);
ha ha4(p[160], s[13], s[14], c[14]);

fa fa10(p[6], p[37], c[10], s[15], c[15]);
fa fa11(p[68], s[15], c[11], s[16], c[16]);
fa fa12(p[99], s[16], c[12], s[17], c[17]);
fa fa13(p[130], s[17], c[13], s[18], c[18]);
fa fa14(p[161], s[18], c[14], s[19], c[19]);
ha ha5(p[192], s[19], s[20], c[20]);

fa fa15(p[7], p[38], c[15], s[21], c[21]);
fa fa16(p[69], s[21], c[16], s[22], c[22]);
fa fa17(p[100], s[22], c[17], s[23], c[23]);
fa fa18(p[131], s[23], c[18], s[24], c[24]);
fa fa19(p[162], s[24], c[19], s[25], c[25]);
fa fa20(p[193], s[25], c[20], s[26], c[26]);
ha ha6(p[224], s[26], s[27], c[27]);

fa fa21(p[8], p[39], c[21], s[28], c[28]);
fa fa22(p[70], s[28], c[22], s[29], c[29]);
fa fa23(p[101], s[29], c[23], s[30], c[30]);
fa fa24(p[132], s[30], c[24], s[31], c[31]);
fa fa25(p[163], s[31], c[25], s[32], c[32]);
fa fa26(p[194], s[32], c[26], s[33], c[33]);
fa fa27(p[225], s[33], c[27], s[34], c[34]);
ha ha7(p[256], s[34], s[35], c[35]);

fa fa28(p[9], p[40], c[28], s[36], c[36]);
fa fa29(p[71], s[36], c[29], s[37], c[37]);
fa fa30(p[102], s[37], c[30], s[38], c[38]);
fa fa31(p[133], s[38], c[31], s[39], c[39]);
fa fa32(p[164], s[39], c[32], s[40], c[40]);
fa fa33(p[195], s[40], c[33], s[41], c[41]);
fa fa34(p[226], s[41], c[34], s[42], c[42]);
fa fa35(p[257], s[42], c[35], s[43], c[43]);
ha ha8(p[288], s[43], s[44], c[44]);

fa fa36(p[10], p[41], c[36], s[45], c[45]);
fa fa37(p[72], s[45], c[37], s[46], c[46]);
fa fa38(p[103], s[46], c[38], s[47], c[47]);
fa fa39(p[134], s[47], c[39], s[48], c[48]);
fa fa40(p[165], s[48], c[40], s[49], c[49]);
fa fa41(p[196], s[49], c[41], s[50], c[50]);
fa fa42(p[227], s[50], c[42], s[51], c[51]);
fa fa43(p[258], s[51], c[43], s[52], c[52]);
fa fa44(p[289], s[52], c[44], s[53], c[53]);
ha ha9(p[320], s[53], s[54], c[54]);

fa fa45(p[11], p[42], c[45], s[55], c[55]);
fa fa46(p[73], s[55], c[46], s[56], c[56]);
fa fa47(p[104], s[56], c[47], s[57], c[57]);
fa fa48(p[135], s[57], c[48], s[58], c[58]);
fa fa49(p[166], s[58], c[49], s[59], c[59]);
fa fa50(p[197], s[59], c[50], s[60], c[60]);
fa fa51(p[228], s[60], c[51], s[61], c[61]);
fa fa52(p[259], s[61], c[52], s[62], c[62]);
fa fa53(p[290], s[62], c[53], s[63], c[63]);
fa fa54(p[321], s[63], c[54], s[64], c[64]);
ha ha10(p[352], s[64], s[65], c[65]);

fa fa55(p[12], p[43], c[55], s[66], c[66]);
fa fa56(p[74], s[66], c[56], s[67], c[67]);
fa fa57(p[105], s[67], c[57], s[68], c[68]);
fa fa58(p[136], s[68], c[58], s[69], c[69]);
fa fa59(p[167], s[69], c[59], s[70], c[70]);
fa fa60(p[198], s[70], c[60], s[71], c[71]);
fa fa61(p[229], s[71], c[61], s[72], c[72]);
fa fa62(p[260], s[72], c[62], s[73], c[73]);
fa fa63(p[291], s[73], c[63], s[74], c[74]);
fa fa64(p[322], s[74], c[64], s[75], c[75]);
fa fa65(p[353], s[75], c[65], s[76], c[76]);
ha ha11(p[384], s[76], s[77], c[77]);

fa fa66(p[13], p[44], c[66], s[78], c[78]);
fa fa67(p[75], s[78], c[67], s[79], c[79]);
fa fa68(p[106], s[79], c[68], s[80], c[80]);
fa fa69(p[137], s[80], c[69], s[81], c[81]);
fa fa70(p[168], s[81], c[70], s[82], c[82]);
fa fa71(p[199], s[82], c[71], s[83], c[83]);
fa fa72(p[230], s[83], c[72], s[84], c[84]);
fa fa73(p[261], s[84], c[73], s[85], c[85]);
fa fa74(p[292], s[85], c[74], s[86], c[86]);
fa fa75(p[323], s[86], c[75], s[87], c[87]);
fa fa76(p[354], s[87], c[76], s[88], c[88]);
fa fa77(p[385], s[88], c[77], s[89], c[89]);
ha ha12(p[416], s[89], s[90], c[90]);

fa fa78(p[14], p[45], c[78], s[91], c[91]);
fa fa79(p[76], s[91], c[79], s[92], c[92]);
fa fa80(p[107], s[92], c[80], s[93], c[93]);
fa fa81(p[138], s[93], c[81], s[94], c[94]);
fa fa82(p[169], s[94], c[82], s[95], c[95]);
fa fa83(p[200], s[95], c[83], s[96], c[96]);
fa fa84(p[231], s[96], c[84], s[97], c[97]);
fa fa85(p[262], s[97], c[85], s[98], c[98]);
fa fa86(p[293], s[98], c[86], s[99], c[99]);
fa fa87(p[324], s[99], c[87], s[100], c[100]);
fa fa88(p[355], s[100], c[88], s[101], c[101]);
fa fa89(p[386], s[101], c[89], s[102], c[102]);
fa fa90(p[417], s[102], c[90], s[103], c[103]);
ha ha13(p[448], s[103], s[104], c[104]);

fa fa91(p[15], p[46], c[91], s[105], c[105]);
fa fa92(p[77], s[105], c[92], s[106], c[106]);
fa fa93(p[108], s[106], c[93], s[107], c[107]);
fa fa94(p[139], s[107], c[94], s[108], c[108]);
fa fa95(p[170], s[108], c[95], s[109], c[109]);
fa fa96(p[201], s[109], c[96], s[110], c[110]);
fa fa97(p[232], s[110], c[97], s[111], c[111]);
fa fa98(p[263], s[111], c[98], s[112], c[112]);
fa fa99(p[294], s[112], c[99], s[113], c[113]);
fa fa100(p[325], s[113], c[100], s[114], c[114]);
fa fa101(p[356], s[114], c[101], s[115], c[115]);
fa fa102(p[387], s[115], c[102], s[116], c[116]);
fa fa103(p[418], s[116], c[103], s[117], c[117]);
fa fa104(p[449], s[117], c[104], s[118], c[118]);
ha ha14(p[480], s[118], s[119], c[119]);

fa fa105(p[16], p[47], c[105], s[120], c[120]);
fa fa106(p[78], s[120], c[106], s[121], c[121]);
fa fa107(p[109], s[121], c[107], s[122], c[122]);
fa fa108(p[140], s[122], c[108], s[123], c[123]);
fa fa109(p[171], s[123], c[109], s[124], c[124]);
fa fa110(p[202], s[124], c[110], s[125], c[125]);
fa fa111(p[233], s[125], c[111], s[126], c[126]);
fa fa112(p[264], s[126], c[112], s[127], c[127]);
fa fa113(p[295], s[127], c[113], s[128], c[128]);
fa fa114(p[326], s[128], c[114], s[129], c[129]);
fa fa115(p[357], s[129], c[115], s[130], c[130]);
fa fa116(p[388], s[130], c[116], s[131], c[131]);
fa fa117(p[419], s[131], c[117], s[132], c[132]);
fa fa118(p[450], s[132], c[118], s[133], c[133]);
fa fa119(p[481], s[133], c[119], s[134], c[134]);
ha ha15(p[512], s[134], s[135], c[135]);

fa fa120(p[17], p[48], c[120], s[136], c[136]);
fa fa121(p[79], s[136], c[121], s[137], c[137]);
fa fa122(p[110], s[137], c[122], s[138], c[138]);
fa fa123(p[141], s[138], c[123], s[139], c[139]);
fa fa124(p[172], s[139], c[124], s[140], c[140]);
fa fa125(p[203], s[140], c[125], s[141], c[141]);
fa fa126(p[234], s[141], c[126], s[142], c[142]);
fa fa127(p[265], s[142], c[127], s[143], c[143]);
fa fa128(p[296], s[143], c[128], s[144], c[144]);
fa fa129(p[327], s[144], c[129], s[145], c[145]);
fa fa130(p[358], s[145], c[130], s[146], c[146]);
fa fa131(p[389], s[146], c[131], s[147], c[147]);
fa fa132(p[420], s[147], c[132], s[148], c[148]);
fa fa133(p[451], s[148], c[133], s[149], c[149]);
fa fa134(p[482], s[149], c[134], s[150], c[150]);
fa fa135(p[513], s[150], c[135], s[151], c[151]);
ha ha16(p[544], s[151], s[152], c[152]);

fa fa136(p[18], p[49], c[136], s[153], c[153]);
fa fa137(p[80], s[153], c[137], s[154], c[154]);
fa fa138(p[111], s[154], c[138], s[155], c[155]);
fa fa139(p[142], s[155], c[139], s[156], c[156]);
fa fa140(p[173], s[156], c[140], s[157], c[157]);
fa fa141(p[204], s[157], c[141], s[158], c[158]);
fa fa142(p[235], s[158], c[142], s[159], c[159]);
fa fa143(p[266], s[159], c[143], s[160], c[160]);
fa fa144(p[297], s[160], c[144], s[161], c[161]);
fa fa145(p[328], s[161], c[145], s[162], c[162]);
fa fa146(p[359], s[162], c[146], s[163], c[163]);
fa fa147(p[390], s[163], c[147], s[164], c[164]);
fa fa148(p[421], s[164], c[148], s[165], c[165]);
fa fa149(p[452], s[165], c[149], s[166], c[166]);
fa fa150(p[483], s[166], c[150], s[167], c[167]);
fa fa151(p[514], s[167], c[151], s[168], c[168]);
fa fa152(p[545], s[168], c[152], s[169], c[169]);
ha ha17(p[576], s[169], s[170], c[170]);

fa fa153(p[19], p[50], c[153], s[171], c[171]);
fa fa154(p[81], s[171], c[154], s[172], c[172]);
fa fa155(p[112], s[172], c[155], s[173], c[173]);
fa fa156(p[143], s[173], c[156], s[174], c[174]);
fa fa157(p[174], s[174], c[157], s[175], c[175]);
fa fa158(p[205], s[175], c[158], s[176], c[176]);
fa fa159(p[236], s[176], c[159], s[177], c[177]);
fa fa160(p[267], s[177], c[160], s[178], c[178]);
fa fa161(p[298], s[178], c[161], s[179], c[179]);
fa fa162(p[329], s[179], c[162], s[180], c[180]);
fa fa163(p[360], s[180], c[163], s[181], c[181]);
fa fa164(p[391], s[181], c[164], s[182], c[182]);
fa fa165(p[422], s[182], c[165], s[183], c[183]);
fa fa166(p[453], s[183], c[166], s[184], c[184]);
fa fa167(p[484], s[184], c[167], s[185], c[185]);
fa fa168(p[515], s[185], c[168], s[186], c[186]);
fa fa169(p[546], s[186], c[169], s[187], c[187]);
fa fa170(p[577], s[187], c[170], s[188], c[188]);
ha ha18(p[608], s[188], s[189], c[189]);

fa fa171(p[20], p[51], c[171], s[190], c[190]);
fa fa172(p[82], s[190], c[172], s[191], c[191]);
fa fa173(p[113], s[191], c[173], s[192], c[192]);
fa fa174(p[144], s[192], c[174], s[193], c[193]);
fa fa175(p[175], s[193], c[175], s[194], c[194]);
fa fa176(p[206], s[194], c[176], s[195], c[195]);
fa fa177(p[237], s[195], c[177], s[196], c[196]);
fa fa178(p[268], s[196], c[178], s[197], c[197]);
fa fa179(p[299], s[197], c[179], s[198], c[198]);
fa fa180(p[330], s[198], c[180], s[199], c[199]);
fa fa181(p[361], s[199], c[181], s[200], c[200]);
fa fa182(p[392], s[200], c[182], s[201], c[201]);
fa fa183(p[423], s[201], c[183], s[202], c[202]);
fa fa184(p[454], s[202], c[184], s[203], c[203]);
fa fa185(p[485], s[203], c[185], s[204], c[204]);
fa fa186(p[516], s[204], c[186], s[205], c[205]);
fa fa187(p[547], s[205], c[187], s[206], c[206]);
fa fa188(p[578], s[206], c[188], s[207], c[207]);
fa fa189(p[609], s[207], c[189], s[208], c[208]);
ha ha19(p[640], s[208], s[209], c[209]);

fa fa190(p[21], p[52], c[190], s[210], c[210]);
fa fa191(p[83], s[210], c[191], s[211], c[211]);
fa fa192(p[114], s[211], c[192], s[212], c[212]);
fa fa193(p[145], s[212], c[193], s[213], c[213]);
fa fa194(p[176], s[213], c[194], s[214], c[214]);
fa fa195(p[207], s[214], c[195], s[215], c[215]);
fa fa196(p[238], s[215], c[196], s[216], c[216]);
fa fa197(p[269], s[216], c[197], s[217], c[217]);
fa fa198(p[300], s[217], c[198], s[218], c[218]);
fa fa199(p[331], s[218], c[199], s[219], c[219]);
fa fa200(p[362], s[219], c[200], s[220], c[220]);
fa fa201(p[393], s[220], c[201], s[221], c[221]);
fa fa202(p[424], s[221], c[202], s[222], c[222]);
fa fa203(p[455], s[222], c[203], s[223], c[223]);
fa fa204(p[486], s[223], c[204], s[224], c[224]);
fa fa205(p[517], s[224], c[205], s[225], c[225]);
fa fa206(p[548], s[225], c[206], s[226], c[226]);
fa fa207(p[579], s[226], c[207], s[227], c[227]);
fa fa208(p[610], s[227], c[208], s[228], c[228]);
fa fa209(p[641], s[228], c[209], s[229], c[229]);
ha ha20(p[672], s[229], s[230], c[230]);

fa fa210(p[22], p[53], c[210], s[231], c[231]);
fa fa211(p[84], s[231], c[211], s[232], c[232]);
fa fa212(p[115], s[232], c[212], s[233], c[233]);
fa fa213(p[146], s[233], c[213], s[234], c[234]);
fa fa214(p[177], s[234], c[214], s[235], c[235]);
fa fa215(p[208], s[235], c[215], s[236], c[236]);
fa fa216(p[239], s[236], c[216], s[237], c[237]);
fa fa217(p[270], s[237], c[217], s[238], c[238]);
fa fa218(p[301], s[238], c[218], s[239], c[239]);
fa fa219(p[332], s[239], c[219], s[240], c[240]);
fa fa220(p[363], s[240], c[220], s[241], c[241]);
fa fa221(p[394], s[241], c[221], s[242], c[242]);
fa fa222(p[425], s[242], c[222], s[243], c[243]);
fa fa223(p[456], s[243], c[223], s[244], c[244]);
fa fa224(p[487], s[244], c[224], s[245], c[245]);
fa fa225(p[518], s[245], c[225], s[246], c[246]);
fa fa226(p[549], s[246], c[226], s[247], c[247]);
fa fa227(p[580], s[247], c[227], s[248], c[248]);
fa fa228(p[611], s[248], c[228], s[249], c[249]);
fa fa229(p[642], s[249], c[229], s[250], c[250]);
fa fa230(p[673], s[250], c[230], s[251], c[251]);
ha ha21(p[704], s[251], s[252], c[252]);

fa fa231(p[23], p[54], c[231], s[253], c[253]);
fa fa232(p[85], s[253], c[232], s[254], c[254]);
fa fa233(p[116], s[254], c[233], s[255], c[255]);
fa fa234(p[147], s[255], c[234], s[256], c[256]);
fa fa235(p[178], s[256], c[235], s[257], c[257]);
fa fa236(p[209], s[257], c[236], s[258], c[258]);
fa fa237(p[240], s[258], c[237], s[259], c[259]);
fa fa238(p[271], s[259], c[238], s[260], c[260]);
fa fa239(p[302], s[260], c[239], s[261], c[261]);
fa fa240(p[333], s[261], c[240], s[262], c[262]);
fa fa241(p[364], s[262], c[241], s[263], c[263]);
fa fa242(p[395], s[263], c[242], s[264], c[264]);
fa fa243(p[426], s[264], c[243], s[265], c[265]);
fa fa244(p[457], s[265], c[244], s[266], c[266]);
fa fa245(p[488], s[266], c[245], s[267], c[267]);
fa fa246(p[519], s[267], c[246], s[268], c[268]);
fa fa247(p[550], s[268], c[247], s[269], c[269]);
fa fa248(p[581], s[269], c[248], s[270], c[270]);
fa fa249(p[612], s[270], c[249], s[271], c[271]);
fa fa250(p[643], s[271], c[250], s[272], c[272]);
fa fa251(p[674], s[272], c[251], s[273], c[273]);
fa fa252(p[705], s[273], c[252], s[274], c[274]);
ha ha22(p[736], s[274], s[275], c[275]);

fa fa253(p[24], p[55], c[253], s[276], c[276]);
fa fa254(p[86], s[276], c[254], s[277], c[277]);
fa fa255(p[117], s[277], c[255], s[278], c[278]);
fa fa256(p[148], s[278], c[256], s[279], c[279]);
fa fa257(p[179], s[279], c[257], s[280], c[280]);
fa fa258(p[210], s[280], c[258], s[281], c[281]);
fa fa259(p[241], s[281], c[259], s[282], c[282]);
fa fa260(p[272], s[282], c[260], s[283], c[283]);
fa fa261(p[303], s[283], c[261], s[284], c[284]);
fa fa262(p[334], s[284], c[262], s[285], c[285]);
fa fa263(p[365], s[285], c[263], s[286], c[286]);
fa fa264(p[396], s[286], c[264], s[287], c[287]);
fa fa265(p[427], s[287], c[265], s[288], c[288]);
fa fa266(p[458], s[288], c[266], s[289], c[289]);
fa fa267(p[489], s[289], c[267], s[290], c[290]);
fa fa268(p[520], s[290], c[268], s[291], c[291]);
fa fa269(p[551], s[291], c[269], s[292], c[292]);
fa fa270(p[582], s[292], c[270], s[293], c[293]);
fa fa271(p[613], s[293], c[271], s[294], c[294]);
fa fa272(p[644], s[294], c[272], s[295], c[295]);
fa fa273(p[675], s[295], c[273], s[296], c[296]);
fa fa274(p[706], s[296], c[274], s[297], c[297]);
fa fa275(p[737], s[297], c[275], s[298], c[298]);
ha ha23(p[768], s[298], s[299], c[299]);

fa fa276(p[25], p[56], c[276], s[300], c[300]);
fa fa277(p[87], s[300], c[277], s[301], c[301]);
fa fa278(p[118], s[301], c[278], s[302], c[302]);
fa fa279(p[149], s[302], c[279], s[303], c[303]);
fa fa280(p[180], s[303], c[280], s[304], c[304]);
fa fa281(p[211], s[304], c[281], s[305], c[305]);
fa fa282(p[242], s[305], c[282], s[306], c[306]);
fa fa283(p[273], s[306], c[283], s[307], c[307]);
fa fa284(p[304], s[307], c[284], s[308], c[308]);
fa fa285(p[335], s[308], c[285], s[309], c[309]);
fa fa286(p[366], s[309], c[286], s[310], c[310]);
fa fa287(p[397], s[310], c[287], s[311], c[311]);
fa fa288(p[428], s[311], c[288], s[312], c[312]);
fa fa289(p[459], s[312], c[289], s[313], c[313]);
fa fa290(p[490], s[313], c[290], s[314], c[314]);
fa fa291(p[521], s[314], c[291], s[315], c[315]);
fa fa292(p[552], s[315], c[292], s[316], c[316]);
fa fa293(p[583], s[316], c[293], s[317], c[317]);
fa fa294(p[614], s[317], c[294], s[318], c[318]);
fa fa295(p[645], s[318], c[295], s[319], c[319]);
fa fa296(p[676], s[319], c[296], s[320], c[320]);
fa fa297(p[707], s[320], c[297], s[321], c[321]);
fa fa298(p[738], s[321], c[298], s[322], c[322]);
fa fa299(p[769], s[322], c[299], s[323], c[323]);
ha ha24(p[800], s[323], s[324], c[324]);

fa fa300(p[26], p[57], c[300], s[325], c[325]);
fa fa301(p[88], s[325], c[301], s[326], c[326]);
fa fa302(p[119], s[326], c[302], s[327], c[327]);
fa fa303(p[150], s[327], c[303], s[328], c[328]);
fa fa304(p[181], s[328], c[304], s[329], c[329]);
fa fa305(p[212], s[329], c[305], s[330], c[330]);
fa fa306(p[243], s[330], c[306], s[331], c[331]);
fa fa307(p[274], s[331], c[307], s[332], c[332]);
fa fa308(p[305], s[332], c[308], s[333], c[333]);
fa fa309(p[336], s[333], c[309], s[334], c[334]);
fa fa310(p[367], s[334], c[310], s[335], c[335]);
fa fa311(p[398], s[335], c[311], s[336], c[336]);
fa fa312(p[429], s[336], c[312], s[337], c[337]);
fa fa313(p[460], s[337], c[313], s[338], c[338]);
fa fa314(p[491], s[338], c[314], s[339], c[339]);
fa fa315(p[522], s[339], c[315], s[340], c[340]);
fa fa316(p[553], s[340], c[316], s[341], c[341]);
fa fa317(p[584], s[341], c[317], s[342], c[342]);
fa fa318(p[615], s[342], c[318], s[343], c[343]);
fa fa319(p[646], s[343], c[319], s[344], c[344]);
fa fa320(p[677], s[344], c[320], s[345], c[345]);
fa fa321(p[708], s[345], c[321], s[346], c[346]);
fa fa322(p[739], s[346], c[322], s[347], c[347]);
fa fa323(p[770], s[347], c[323], s[348], c[348]);
fa fa324(p[801], s[348], c[324], s[349], c[349]);
ha ha25(p[832], s[349], s[350], c[350]);

fa fa325(p[27], p[58], c[325], s[351], c[351]);
fa fa326(p[89], s[351], c[326], s[352], c[352]);
fa fa327(p[120], s[352], c[327], s[353], c[353]);
fa fa328(p[151], s[353], c[328], s[354], c[354]);
fa fa329(p[182], s[354], c[329], s[355], c[355]);
fa fa330(p[213], s[355], c[330], s[356], c[356]);
fa fa331(p[244], s[356], c[331], s[357], c[357]);
fa fa332(p[275], s[357], c[332], s[358], c[358]);
fa fa333(p[306], s[358], c[333], s[359], c[359]);
fa fa334(p[337], s[359], c[334], s[360], c[360]);
fa fa335(p[368], s[360], c[335], s[361], c[361]);
fa fa336(p[399], s[361], c[336], s[362], c[362]);
fa fa337(p[430], s[362], c[337], s[363], c[363]);
fa fa338(p[461], s[363], c[338], s[364], c[364]);
fa fa339(p[492], s[364], c[339], s[365], c[365]);
fa fa340(p[523], s[365], c[340], s[366], c[366]);
fa fa341(p[554], s[366], c[341], s[367], c[367]);
fa fa342(p[585], s[367], c[342], s[368], c[368]);
fa fa343(p[616], s[368], c[343], s[369], c[369]);
fa fa344(p[647], s[369], c[344], s[370], c[370]);
fa fa345(p[678], s[370], c[345], s[371], c[371]);
fa fa346(p[709], s[371], c[346], s[372], c[372]);
fa fa347(p[740], s[372], c[347], s[373], c[373]);
fa fa348(p[771], s[373], c[348], s[374], c[374]);
fa fa349(p[802], s[374], c[349], s[375], c[375]);
fa fa350(p[833], s[375], c[350], s[376], c[376]);
ha ha26(p[864], s[376], s[377], c[377]);

fa fa351(p[28], p[59], c[351], s[378], c[378]);
fa fa352(p[90], s[378], c[352], s[379], c[379]);
fa fa353(p[121], s[379], c[353], s[380], c[380]);
fa fa354(p[152], s[380], c[354], s[381], c[381]);
fa fa355(p[183], s[381], c[355], s[382], c[382]);
fa fa356(p[214], s[382], c[356], s[383], c[383]);
fa fa357(p[245], s[383], c[357], s[384], c[384]);
fa fa358(p[276], s[384], c[358], s[385], c[385]);
fa fa359(p[307], s[385], c[359], s[386], c[386]);
fa fa360(p[338], s[386], c[360], s[387], c[387]);
fa fa361(p[369], s[387], c[361], s[388], c[388]);
fa fa362(p[400], s[388], c[362], s[389], c[389]);
fa fa363(p[431], s[389], c[363], s[390], c[390]);
fa fa364(p[462], s[390], c[364], s[391], c[391]);
fa fa365(p[493], s[391], c[365], s[392], c[392]);
fa fa366(p[524], s[392], c[366], s[393], c[393]);
fa fa367(p[555], s[393], c[367], s[394], c[394]);
fa fa368(p[586], s[394], c[368], s[395], c[395]);
fa fa369(p[617], s[395], c[369], s[396], c[396]);
fa fa370(p[648], s[396], c[370], s[397], c[397]);
fa fa371(p[679], s[397], c[371], s[398], c[398]);
fa fa372(p[710], s[398], c[372], s[399], c[399]);
fa fa373(p[741], s[399], c[373], s[400], c[400]);
fa fa374(p[772], s[400], c[374], s[401], c[401]);
fa fa375(p[803], s[401], c[375], s[402], c[402]);
fa fa376(p[834], s[402], c[376], s[403], c[403]);
fa fa377(p[865], s[403], c[377], s[404], c[404]);
ha ha27(p[896], s[404], s[405], c[405]);

fa fa378(p[29], p[60], c[378], s[406], c[406]);
fa fa379(p[91], s[406], c[379], s[407], c[407]);
fa fa380(p[122], s[407], c[380], s[408], c[408]);
fa fa381(p[153], s[408], c[381], s[409], c[409]);
fa fa382(p[184], s[409], c[382], s[410], c[410]);
fa fa383(p[215], s[410], c[383], s[411], c[411]);
fa fa384(p[246], s[411], c[384], s[412], c[412]);
fa fa385(p[277], s[412], c[385], s[413], c[413]);
fa fa386(p[308], s[413], c[386], s[414], c[414]);
fa fa387(p[339], s[414], c[387], s[415], c[415]);
fa fa388(p[370], s[415], c[388], s[416], c[416]);
fa fa389(p[401], s[416], c[389], s[417], c[417]);
fa fa390(p[432], s[417], c[390], s[418], c[418]);
fa fa391(p[463], s[418], c[391], s[419], c[419]);
fa fa392(p[494], s[419], c[392], s[420], c[420]);
fa fa393(p[525], s[420], c[393], s[421], c[421]);
fa fa394(p[556], s[421], c[394], s[422], c[422]);
fa fa395(p[587], s[422], c[395], s[423], c[423]);
fa fa396(p[618], s[423], c[396], s[424], c[424]);
fa fa397(p[649], s[424], c[397], s[425], c[425]);
fa fa398(p[680], s[425], c[398], s[426], c[426]);
fa fa399(p[711], s[426], c[399], s[427], c[427]);
fa fa400(p[742], s[427], c[400], s[428], c[428]);
fa fa401(p[773], s[428], c[401], s[429], c[429]);
fa fa402(p[804], s[429], c[402], s[430], c[430]);
fa fa403(p[835], s[430], c[403], s[431], c[431]);
fa fa404(p[866], s[431], c[404], s[432], c[432]);
fa fa405(p[897], s[432], c[405], s[433], c[433]);
ha ha28(p[928], s[433], s[434], c[434]);

fa fa406(p[30], p[61], c[406], s[435], c[435]);
fa fa407(p[92], s[435], c[407], s[436], c[436]);
fa fa408(p[123], s[436], c[408], s[437], c[437]);
fa fa409(p[154], s[437], c[409], s[438], c[438]);
fa fa410(p[185], s[438], c[410], s[439], c[439]);
fa fa411(p[216], s[439], c[411], s[440], c[440]);
fa fa412(p[247], s[440], c[412], s[441], c[441]);
fa fa413(p[278], s[441], c[413], s[442], c[442]);
fa fa414(p[309], s[442], c[414], s[443], c[443]);
fa fa415(p[340], s[443], c[415], s[444], c[444]);
fa fa416(p[371], s[444], c[416], s[445], c[445]);
fa fa417(p[402], s[445], c[417], s[446], c[446]);
fa fa418(p[433], s[446], c[418], s[447], c[447]);
fa fa419(p[464], s[447], c[419], s[448], c[448]);
fa fa420(p[495], s[448], c[420], s[449], c[449]);
fa fa421(p[526], s[449], c[421], s[450], c[450]);
fa fa422(p[557], s[450], c[422], s[451], c[451]);
fa fa423(p[588], s[451], c[423], s[452], c[452]);
fa fa424(p[619], s[452], c[424], s[453], c[453]);
fa fa425(p[650], s[453], c[425], s[454], c[454]);
fa fa426(p[681], s[454], c[426], s[455], c[455]);
fa fa427(p[712], s[455], c[427], s[456], c[456]);
fa fa428(p[743], s[456], c[428], s[457], c[457]);
fa fa429(p[774], s[457], c[429], s[458], c[458]);
fa fa430(p[805], s[458], c[430], s[459], c[459]);
fa fa431(p[836], s[459], c[431], s[460], c[460]);
fa fa432(p[867], s[460], c[432], s[461], c[461]);
fa fa433(p[898], s[461], c[433], s[462], c[462]);
fa fa434(p[929], s[462], c[434], s[463], c[463]);
ha ha29(p[960], s[463], s[464], c[464]);

fa fa435(p[31], p[62], c[435], s[465], c[465]);
fa fa436(p[93], s[465], c[436], s[466], c[466]);
fa fa437(p[124], s[466], c[437], s[467], c[467]);
fa fa438(p[155], s[467], c[438], s[468], c[468]);
fa fa439(p[186], s[468], c[439], s[469], c[469]);
fa fa440(p[217], s[469], c[440], s[470], c[470]);
fa fa441(p[248], s[470], c[441], s[471], c[471]);
fa fa442(p[279], s[471], c[442], s[472], c[472]);
fa fa443(p[310], s[472], c[443], s[473], c[473]);
fa fa444(p[341], s[473], c[444], s[474], c[474]);
fa fa445(p[372], s[474], c[445], s[475], c[475]);
fa fa446(p[403], s[475], c[446], s[476], c[476]);
fa fa447(p[434], s[476], c[447], s[477], c[477]);
fa fa448(p[465], s[477], c[448], s[478], c[478]);
fa fa449(p[496], s[478], c[449], s[479], c[479]);
fa fa450(p[527], s[479], c[450], s[480], c[480]);
fa fa451(p[558], s[480], c[451], s[481], c[481]);
fa fa452(p[589], s[481], c[452], s[482], c[482]);
fa fa453(p[620], s[482], c[453], s[483], c[483]);
fa fa454(p[651], s[483], c[454], s[484], c[484]);
fa fa455(p[682], s[484], c[455], s[485], c[485]);
fa fa456(p[713], s[485], c[456], s[486], c[486]);
fa fa457(p[744], s[486], c[457], s[487], c[487]);
fa fa458(p[775], s[487], c[458], s[488], c[488]);
fa fa459(p[806], s[488], c[459], s[489], c[489]);
fa fa460(p[837], s[489], c[460], s[490], c[490]);
fa fa461(p[868], s[490], c[461], s[491], c[491]);
fa fa462(p[899], s[491], c[462], s[492], c[492]);
fa fa463(p[930], s[492], c[463], s[493], c[493]);
fa fa464(p[961], s[493], c[464], s[494], c[494]);
ha ha30(p[992], s[494], s[495], c[495]);

fa fa465(p[63], c[465], c[466], s[496], c[496]);
fa fa466(p[94], s[496], c[467], s[497], c[497]);
fa fa467(p[125], s[497], c[468], s[498], c[498]);
fa fa468(p[156], s[498], c[469], s[499], c[499]);
fa fa469(p[187], s[499], c[470], s[500], c[500]);
fa fa470(p[218], s[500], c[471], s[501], c[501]);
fa fa471(p[249], s[501], c[472], s[502], c[502]);
fa fa472(p[280], s[502], c[473], s[503], c[503]);
fa fa473(p[311], s[503], c[474], s[504], c[504]);
fa fa474(p[342], s[504], c[475], s[505], c[505]);
fa fa475(p[373], s[505], c[476], s[506], c[506]);
fa fa476(p[404], s[506], c[477], s[507], c[507]);
fa fa477(p[435], s[507], c[478], s[508], c[508]);
fa fa478(p[466], s[508], c[479], s[509], c[509]);
fa fa479(p[497], s[509], c[480], s[510], c[510]);
fa fa480(p[528], s[510], c[481], s[511], c[511]);
fa fa481(p[559], s[511], c[482], s[512], c[512]);
fa fa482(p[590], s[512], c[483], s[513], c[513]);
fa fa483(p[621], s[513], c[484], s[514], c[514]);
fa fa484(p[652], s[514], c[485], s[515], c[515]);
fa fa485(p[683], s[515], c[486], s[516], c[516]);
fa fa486(p[714], s[516], c[487], s[517], c[517]);
fa fa487(p[745], s[517], c[488], s[518], c[518]);
fa fa488(p[776], s[518], c[489], s[519], c[519]);
fa fa489(p[807], s[519], c[490], s[520], c[520]);
fa fa490(p[838], s[520], c[491], s[521], c[521]);
fa fa491(p[869], s[521], c[492], s[522], c[522]);
fa fa492(p[900], s[522], c[493], s[523], c[523]);
fa fa493(p[931], s[523], c[494], s[524], c[524]);
fa fa494(p[962], s[524], c[495], s[525], c[525]);
ha ha31(p[993], s[525], s[526], c[526]);

fa fa495(p[95], c[496], c[497], s[527], c[527]);
fa fa496(p[126], s[527], c[498], s[528], c[528]);
fa fa497(p[157], s[528], c[499], s[529], c[529]);
fa fa498(p[188], s[529], c[500], s[530], c[530]);
fa fa499(p[219], s[530], c[501], s[531], c[531]);
fa fa500(p[250], s[531], c[502], s[532], c[532]);
fa fa501(p[281], s[532], c[503], s[533], c[533]);
fa fa502(p[312], s[533], c[504], s[534], c[534]);
fa fa503(p[343], s[534], c[505], s[535], c[535]);
fa fa504(p[374], s[535], c[506], s[536], c[536]);
fa fa505(p[405], s[536], c[507], s[537], c[537]);
fa fa506(p[436], s[537], c[508], s[538], c[538]);
fa fa507(p[467], s[538], c[509], s[539], c[539]);
fa fa508(p[498], s[539], c[510], s[540], c[540]);
fa fa509(p[529], s[540], c[511], s[541], c[541]);
fa fa510(p[560], s[541], c[512], s[542], c[542]);
fa fa511(p[591], s[542], c[513], s[543], c[543]);
fa fa512(p[622], s[543], c[514], s[544], c[544]);
fa fa513(p[653], s[544], c[515], s[545], c[545]);
fa fa514(p[684], s[545], c[516], s[546], c[546]);
fa fa515(p[715], s[546], c[517], s[547], c[547]);
fa fa516(p[746], s[547], c[518], s[548], c[548]);
fa fa517(p[777], s[548], c[519], s[549], c[549]);
fa fa518(p[808], s[549], c[520], s[550], c[550]);
fa fa519(p[839], s[550], c[521], s[551], c[551]);
fa fa520(p[870], s[551], c[522], s[552], c[552]);
fa fa521(p[901], s[552], c[523], s[553], c[553]);
fa fa522(p[932], s[553], c[524], s[554], c[554]);
fa fa523(p[963], s[554], c[525], s[555], c[555]);
fa fa524(p[994], s[555], c[526], s[556], c[556]);

fa fa525(p[127], c[527], c[528], s[557], c[557]);
fa fa526(p[158], s[557], c[529], s[558], c[558]);
fa fa527(p[189], s[558], c[530], s[559], c[559]);
fa fa528(p[220], s[559], c[531], s[560], c[560]);
fa fa529(p[251], s[560], c[532], s[561], c[561]);
fa fa530(p[282], s[561], c[533], s[562], c[562]);
fa fa531(p[313], s[562], c[534], s[563], c[563]);
fa fa532(p[344], s[563], c[535], s[564], c[564]);
fa fa533(p[375], s[564], c[536], s[565], c[565]);
fa fa534(p[406], s[565], c[537], s[566], c[566]);
fa fa535(p[437], s[566], c[538], s[567], c[567]);
fa fa536(p[468], s[567], c[539], s[568], c[568]);
fa fa537(p[499], s[568], c[540], s[569], c[569]);
fa fa538(p[530], s[569], c[541], s[570], c[570]);
fa fa539(p[561], s[570], c[542], s[571], c[571]);
fa fa540(p[592], s[571], c[543], s[572], c[572]);
fa fa541(p[623], s[572], c[544], s[573], c[573]);
fa fa542(p[654], s[573], c[545], s[574], c[574]);
fa fa543(p[685], s[574], c[546], s[575], c[575]);
fa fa544(p[716], s[575], c[547], s[576], c[576]);
fa fa545(p[747], s[576], c[548], s[577], c[577]);
fa fa546(p[778], s[577], c[549], s[578], c[578]);
fa fa547(p[809], s[578], c[550], s[579], c[579]);
fa fa548(p[840], s[579], c[551], s[580], c[580]);
fa fa549(p[871], s[580], c[552], s[581], c[581]);
fa fa550(p[902], s[581], c[553], s[582], c[582]);
fa fa551(p[933], s[582], c[554], s[583], c[583]);
fa fa552(p[964], s[583], c[555], s[584], c[584]);
fa fa553(p[995], s[584], c[556], s[585], c[585]);

fa fa554(p[159], c[557], c[558], s[586], c[586]);
fa fa555(p[190], s[586], c[559], s[587], c[587]);
fa fa556(p[221], s[587], c[560], s[588], c[588]);
fa fa557(p[252], s[588], c[561], s[589], c[589]);
fa fa558(p[283], s[589], c[562], s[590], c[590]);
fa fa559(p[314], s[590], c[563], s[591], c[591]);
fa fa560(p[345], s[591], c[564], s[592], c[592]);
fa fa561(p[376], s[592], c[565], s[593], c[593]);
fa fa562(p[407], s[593], c[566], s[594], c[594]);
fa fa563(p[438], s[594], c[567], s[595], c[595]);
fa fa564(p[469], s[595], c[568], s[596], c[596]);
fa fa565(p[500], s[596], c[569], s[597], c[597]);
fa fa566(p[531], s[597], c[570], s[598], c[598]);
fa fa567(p[562], s[598], c[571], s[599], c[599]);
fa fa568(p[593], s[599], c[572], s[600], c[600]);
fa fa569(p[624], s[600], c[573], s[601], c[601]);
fa fa570(p[655], s[601], c[574], s[602], c[602]);
fa fa571(p[686], s[602], c[575], s[603], c[603]);
fa fa572(p[717], s[603], c[576], s[604], c[604]);
fa fa573(p[748], s[604], c[577], s[605], c[605]);
fa fa574(p[779], s[605], c[578], s[606], c[606]);
fa fa575(p[810], s[606], c[579], s[607], c[607]);
fa fa576(p[841], s[607], c[580], s[608], c[608]);
fa fa577(p[872], s[608], c[581], s[609], c[609]);
fa fa578(p[903], s[609], c[582], s[610], c[610]);
fa fa579(p[934], s[610], c[583], s[611], c[611]);
fa fa580(p[965], s[611], c[584], s[612], c[612]);
fa fa581(p[996], s[612], c[585], s[613], c[613]);

fa fa582(p[191], c[586], c[587], s[614], c[614]);
fa fa583(p[222], s[614], c[588], s[615], c[615]);
fa fa584(p[253], s[615], c[589], s[616], c[616]);
fa fa585(p[284], s[616], c[590], s[617], c[617]);
fa fa586(p[315], s[617], c[591], s[618], c[618]);
fa fa587(p[346], s[618], c[592], s[619], c[619]);
fa fa588(p[377], s[619], c[593], s[620], c[620]);
fa fa589(p[408], s[620], c[594], s[621], c[621]);
fa fa590(p[439], s[621], c[595], s[622], c[622]);
fa fa591(p[470], s[622], c[596], s[623], c[623]);
fa fa592(p[501], s[623], c[597], s[624], c[624]);
fa fa593(p[532], s[624], c[598], s[625], c[625]);
fa fa594(p[563], s[625], c[599], s[626], c[626]);
fa fa595(p[594], s[626], c[600], s[627], c[627]);
fa fa596(p[625], s[627], c[601], s[628], c[628]);
fa fa597(p[656], s[628], c[602], s[629], c[629]);
fa fa598(p[687], s[629], c[603], s[630], c[630]);
fa fa599(p[718], s[630], c[604], s[631], c[631]);
fa fa600(p[749], s[631], c[605], s[632], c[632]);
fa fa601(p[780], s[632], c[606], s[633], c[633]);
fa fa602(p[811], s[633], c[607], s[634], c[634]);
fa fa603(p[842], s[634], c[608], s[635], c[635]);
fa fa604(p[873], s[635], c[609], s[636], c[636]);
fa fa605(p[904], s[636], c[610], s[637], c[637]);
fa fa606(p[935], s[637], c[611], s[638], c[638]);
fa fa607(p[966], s[638], c[612], s[639], c[639]);
fa fa608(p[997], s[639], c[613], s[640], c[640]);

fa fa609(p[223], c[614], c[615], s[641], c[641]);
fa fa610(p[254], s[641], c[616], s[642], c[642]);
fa fa611(p[285], s[642], c[617], s[643], c[643]);
fa fa612(p[316], s[643], c[618], s[644], c[644]);
fa fa613(p[347], s[644], c[619], s[645], c[645]);
fa fa614(p[378], s[645], c[620], s[646], c[646]);
fa fa615(p[409], s[646], c[621], s[647], c[647]);
fa fa616(p[440], s[647], c[622], s[648], c[648]);
fa fa617(p[471], s[648], c[623], s[649], c[649]);
fa fa618(p[502], s[649], c[624], s[650], c[650]);
fa fa619(p[533], s[650], c[625], s[651], c[651]);
fa fa620(p[564], s[651], c[626], s[652], c[652]);
fa fa621(p[595], s[652], c[627], s[653], c[653]);
fa fa622(p[626], s[653], c[628], s[654], c[654]);
fa fa623(p[657], s[654], c[629], s[655], c[655]);
fa fa624(p[688], s[655], c[630], s[656], c[656]);
fa fa625(p[719], s[656], c[631], s[657], c[657]);
fa fa626(p[750], s[657], c[632], s[658], c[658]);
fa fa627(p[781], s[658], c[633], s[659], c[659]);
fa fa628(p[812], s[659], c[634], s[660], c[660]);
fa fa629(p[843], s[660], c[635], s[661], c[661]);
fa fa630(p[874], s[661], c[636], s[662], c[662]);
fa fa631(p[905], s[662], c[637], s[663], c[663]);
fa fa632(p[936], s[663], c[638], s[664], c[664]);
fa fa633(p[967], s[664], c[639], s[665], c[665]);
fa fa634(p[998], s[665], c[640], s[666], c[666]);

fa fa635(p[255], c[641], c[642], s[667], c[667]);
fa fa636(p[286], s[667], c[643], s[668], c[668]);
fa fa637(p[317], s[668], c[644], s[669], c[669]);
fa fa638(p[348], s[669], c[645], s[670], c[670]);
fa fa639(p[379], s[670], c[646], s[671], c[671]);
fa fa640(p[410], s[671], c[647], s[672], c[672]);
fa fa641(p[441], s[672], c[648], s[673], c[673]);
fa fa642(p[472], s[673], c[649], s[674], c[674]);
fa fa643(p[503], s[674], c[650], s[675], c[675]);
fa fa644(p[534], s[675], c[651], s[676], c[676]);
fa fa645(p[565], s[676], c[652], s[677], c[677]);
fa fa646(p[596], s[677], c[653], s[678], c[678]);
fa fa647(p[627], s[678], c[654], s[679], c[679]);
fa fa648(p[658], s[679], c[655], s[680], c[680]);
fa fa649(p[689], s[680], c[656], s[681], c[681]);
fa fa650(p[720], s[681], c[657], s[682], c[682]);
fa fa651(p[751], s[682], c[658], s[683], c[683]);
fa fa652(p[782], s[683], c[659], s[684], c[684]);
fa fa653(p[813], s[684], c[660], s[685], c[685]);
fa fa654(p[844], s[685], c[661], s[686], c[686]);
fa fa655(p[875], s[686], c[662], s[687], c[687]);
fa fa656(p[906], s[687], c[663], s[688], c[688]);
fa fa657(p[937], s[688], c[664], s[689], c[689]);
fa fa658(p[968], s[689], c[665], s[690], c[690]);
fa fa659(p[999], s[690], c[666], s[691], c[691]);

fa fa660(p[287], c[667], c[668], s[692], c[692]);
fa fa661(p[318], s[692], c[669], s[693], c[693]);
fa fa662(p[349], s[693], c[670], s[694], c[694]);
fa fa663(p[380], s[694], c[671], s[695], c[695]);
fa fa664(p[411], s[695], c[672], s[696], c[696]);
fa fa665(p[442], s[696], c[673], s[697], c[697]);
fa fa666(p[473], s[697], c[674], s[698], c[698]);
fa fa667(p[504], s[698], c[675], s[699], c[699]);
fa fa668(p[535], s[699], c[676], s[700], c[700]);
fa fa669(p[566], s[700], c[677], s[701], c[701]);
fa fa670(p[597], s[701], c[678], s[702], c[702]);
fa fa671(p[628], s[702], c[679], s[703], c[703]);
fa fa672(p[659], s[703], c[680], s[704], c[704]);
fa fa673(p[690], s[704], c[681], s[705], c[705]);
fa fa674(p[721], s[705], c[682], s[706], c[706]);
fa fa675(p[752], s[706], c[683], s[707], c[707]);
fa fa676(p[783], s[707], c[684], s[708], c[708]);
fa fa677(p[814], s[708], c[685], s[709], c[709]);
fa fa678(p[845], s[709], c[686], s[710], c[710]);
fa fa679(p[876], s[710], c[687], s[711], c[711]);
fa fa680(p[907], s[711], c[688], s[712], c[712]);
fa fa681(p[938], s[712], c[689], s[713], c[713]);
fa fa682(p[969], s[713], c[690], s[714], c[714]);
fa fa683(p[1000], s[714], c[691], s[715], c[715]);

fa fa684(p[319], c[692], c[693], s[716], c[716]);
fa fa685(p[350], s[716], c[694], s[717], c[717]);
fa fa686(p[381], s[717], c[695], s[718], c[718]);
fa fa687(p[412], s[718], c[696], s[719], c[719]);
fa fa688(p[443], s[719], c[697], s[720], c[720]);
fa fa689(p[474], s[720], c[698], s[721], c[721]);
fa fa690(p[505], s[721], c[699], s[722], c[722]);
fa fa691(p[536], s[722], c[700], s[723], c[723]);
fa fa692(p[567], s[723], c[701], s[724], c[724]);
fa fa693(p[598], s[724], c[702], s[725], c[725]);
fa fa694(p[629], s[725], c[703], s[726], c[726]);
fa fa695(p[660], s[726], c[704], s[727], c[727]);
fa fa696(p[691], s[727], c[705], s[728], c[728]);
fa fa697(p[722], s[728], c[706], s[729], c[729]);
fa fa698(p[753], s[729], c[707], s[730], c[730]);
fa fa699(p[784], s[730], c[708], s[731], c[731]);
fa fa700(p[815], s[731], c[709], s[732], c[732]);
fa fa701(p[846], s[732], c[710], s[733], c[733]);
fa fa702(p[877], s[733], c[711], s[734], c[734]);
fa fa703(p[908], s[734], c[712], s[735], c[735]);
fa fa704(p[939], s[735], c[713], s[736], c[736]);
fa fa705(p[970], s[736], c[714], s[737], c[737]);
fa fa706(p[1001], s[737], c[715], s[738], c[738]);

fa fa707(p[351], c[716], c[717], s[739], c[739]);
fa fa708(p[382], s[739], c[718], s[740], c[740]);
fa fa709(p[413], s[740], c[719], s[741], c[741]);
fa fa710(p[444], s[741], c[720], s[742], c[742]);
fa fa711(p[475], s[742], c[721], s[743], c[743]);
fa fa712(p[506], s[743], c[722], s[744], c[744]);
fa fa713(p[537], s[744], c[723], s[745], c[745]);
fa fa714(p[568], s[745], c[724], s[746], c[746]);
fa fa715(p[599], s[746], c[725], s[747], c[747]);
fa fa716(p[630], s[747], c[726], s[748], c[748]);
fa fa717(p[661], s[748], c[727], s[749], c[749]);
fa fa718(p[692], s[749], c[728], s[750], c[750]);
fa fa719(p[723], s[750], c[729], s[751], c[751]);
fa fa720(p[754], s[751], c[730], s[752], c[752]);
fa fa721(p[785], s[752], c[731], s[753], c[753]);
fa fa722(p[816], s[753], c[732], s[754], c[754]);
fa fa723(p[847], s[754], c[733], s[755], c[755]);
fa fa724(p[878], s[755], c[734], s[756], c[756]);
fa fa725(p[909], s[756], c[735], s[757], c[757]);
fa fa726(p[940], s[757], c[736], s[758], c[758]);
fa fa727(p[971], s[758], c[737], s[759], c[759]);
fa fa728(p[1002], s[759], c[738], s[760], c[760]);

fa fa729(p[383], c[739], c[740], s[761], c[761]);
fa fa730(p[414], s[761], c[741], s[762], c[762]);
fa fa731(p[445], s[762], c[742], s[763], c[763]);
fa fa732(p[476], s[763], c[743], s[764], c[764]);
fa fa733(p[507], s[764], c[744], s[765], c[765]);
fa fa734(p[538], s[765], c[745], s[766], c[766]);
fa fa735(p[569], s[766], c[746], s[767], c[767]);
fa fa736(p[600], s[767], c[747], s[768], c[768]);
fa fa737(p[631], s[768], c[748], s[769], c[769]);
fa fa738(p[662], s[769], c[749], s[770], c[770]);
fa fa739(p[693], s[770], c[750], s[771], c[771]);
fa fa740(p[724], s[771], c[751], s[772], c[772]);
fa fa741(p[755], s[772], c[752], s[773], c[773]);
fa fa742(p[786], s[773], c[753], s[774], c[774]);
fa fa743(p[817], s[774], c[754], s[775], c[775]);
fa fa744(p[848], s[775], c[755], s[776], c[776]);
fa fa745(p[879], s[776], c[756], s[777], c[777]);
fa fa746(p[910], s[777], c[757], s[778], c[778]);
fa fa747(p[941], s[778], c[758], s[779], c[779]);
fa fa748(p[972], s[779], c[759], s[780], c[780]);
fa fa749(p[1003], s[780], c[760], s[781], c[781]);

fa fa750(p[415], c[761], c[762], s[782], c[782]);
fa fa751(p[446], s[782], c[763], s[783], c[783]);
fa fa752(p[477], s[783], c[764], s[784], c[784]);
fa fa753(p[508], s[784], c[765], s[785], c[785]);
fa fa754(p[539], s[785], c[766], s[786], c[786]);
fa fa755(p[570], s[786], c[767], s[787], c[787]);
fa fa756(p[601], s[787], c[768], s[788], c[788]);
fa fa757(p[632], s[788], c[769], s[789], c[789]);
fa fa758(p[663], s[789], c[770], s[790], c[790]);
fa fa759(p[694], s[790], c[771], s[791], c[791]);
fa fa760(p[725], s[791], c[772], s[792], c[792]);
fa fa761(p[756], s[792], c[773], s[793], c[793]);
fa fa762(p[787], s[793], c[774], s[794], c[794]);
fa fa763(p[818], s[794], c[775], s[795], c[795]);
fa fa764(p[849], s[795], c[776], s[796], c[796]);
fa fa765(p[880], s[796], c[777], s[797], c[797]);
fa fa766(p[911], s[797], c[778], s[798], c[798]);
fa fa767(p[942], s[798], c[779], s[799], c[799]);
fa fa768(p[973], s[799], c[780], s[800], c[800]);
fa fa769(p[1004], s[800], c[781], s[801], c[801]);

fa fa770(p[447], c[782], c[783], s[802], c[802]);
fa fa771(p[478], s[802], c[784], s[803], c[803]);
fa fa772(p[509], s[803], c[785], s[804], c[804]);
fa fa773(p[540], s[804], c[786], s[805], c[805]);
fa fa774(p[571], s[805], c[787], s[806], c[806]);
fa fa775(p[602], s[806], c[788], s[807], c[807]);
fa fa776(p[633], s[807], c[789], s[808], c[808]);
fa fa777(p[664], s[808], c[790], s[809], c[809]);
fa fa778(p[695], s[809], c[791], s[810], c[810]);
fa fa779(p[726], s[810], c[792], s[811], c[811]);
fa fa780(p[757], s[811], c[793], s[812], c[812]);
fa fa781(p[788], s[812], c[794], s[813], c[813]);
fa fa782(p[819], s[813], c[795], s[814], c[814]);
fa fa783(p[850], s[814], c[796], s[815], c[815]);
fa fa784(p[881], s[815], c[797], s[816], c[816]);
fa fa785(p[912], s[816], c[798], s[817], c[817]);
fa fa786(p[943], s[817], c[799], s[818], c[818]);
fa fa787(p[974], s[818], c[800], s[819], c[819]);
fa fa788(p[1005], s[819], c[801], s[820], c[820]);

fa fa789(p[479], c[802], c[803], s[821], c[821]);
fa fa790(p[510], s[821], c[804], s[822], c[822]);
fa fa791(p[541], s[822], c[805], s[823], c[823]);
fa fa792(p[572], s[823], c[806], s[824], c[824]);
fa fa793(p[603], s[824], c[807], s[825], c[825]);
fa fa794(p[634], s[825], c[808], s[826], c[826]);
fa fa795(p[665], s[826], c[809], s[827], c[827]);
fa fa796(p[696], s[827], c[810], s[828], c[828]);
fa fa797(p[727], s[828], c[811], s[829], c[829]);
fa fa798(p[758], s[829], c[812], s[830], c[830]);
fa fa799(p[789], s[830], c[813], s[831], c[831]);
fa fa800(p[820], s[831], c[814], s[832], c[832]);
fa fa801(p[851], s[832], c[815], s[833], c[833]);
fa fa802(p[882], s[833], c[816], s[834], c[834]);
fa fa803(p[913], s[834], c[817], s[835], c[835]);
fa fa804(p[944], s[835], c[818], s[836], c[836]);
fa fa805(p[975], s[836], c[819], s[837], c[837]);
fa fa806(p[1006], s[837], c[820], s[838], c[838]);

fa fa807(p[511], c[821], c[822], s[839], c[839]);
fa fa808(p[542], s[839], c[823], s[840], c[840]);
fa fa809(p[573], s[840], c[824], s[841], c[841]);
fa fa810(p[604], s[841], c[825], s[842], c[842]);
fa fa811(p[635], s[842], c[826], s[843], c[843]);
fa fa812(p[666], s[843], c[827], s[844], c[844]);
fa fa813(p[697], s[844], c[828], s[845], c[845]);
fa fa814(p[728], s[845], c[829], s[846], c[846]);
fa fa815(p[759], s[846], c[830], s[847], c[847]);
fa fa816(p[790], s[847], c[831], s[848], c[848]);
fa fa817(p[821], s[848], c[832], s[849], c[849]);
fa fa818(p[852], s[849], c[833], s[850], c[850]);
fa fa819(p[883], s[850], c[834], s[851], c[851]);
fa fa820(p[914], s[851], c[835], s[852], c[852]);
fa fa821(p[945], s[852], c[836], s[853], c[853]);
fa fa822(p[976], s[853], c[837], s[854], c[854]);
fa fa823(p[1007], s[854], c[838], s[855], c[855]);

fa fa824(p[543], c[839], c[840], s[856], c[856]);
fa fa825(p[574], s[856], c[841], s[857], c[857]);
fa fa826(p[605], s[857], c[842], s[858], c[858]);
fa fa827(p[636], s[858], c[843], s[859], c[859]);
fa fa828(p[667], s[859], c[844], s[860], c[860]);
fa fa829(p[698], s[860], c[845], s[861], c[861]);
fa fa830(p[729], s[861], c[846], s[862], c[862]);
fa fa831(p[760], s[862], c[847], s[863], c[863]);
fa fa832(p[791], s[863], c[848], s[864], c[864]);
fa fa833(p[822], s[864], c[849], s[865], c[865]);
fa fa834(p[853], s[865], c[850], s[866], c[866]);
fa fa835(p[884], s[866], c[851], s[867], c[867]);
fa fa836(p[915], s[867], c[852], s[868], c[868]);
fa fa837(p[946], s[868], c[853], s[869], c[869]);
fa fa838(p[977], s[869], c[854], s[870], c[870]);
fa fa839(p[1008], s[870], c[855], s[871], c[871]);

fa fa840(p[575], c[856], c[857], s[872], c[872]);
fa fa841(p[606], s[872], c[858], s[873], c[873]);
fa fa842(p[637], s[873], c[859], s[874], c[874]);
fa fa843(p[668], s[874], c[860], s[875], c[875]);
fa fa844(p[699], s[875], c[861], s[876], c[876]);
fa fa845(p[730], s[876], c[862], s[877], c[877]);
fa fa846(p[761], s[877], c[863], s[878], c[878]);
fa fa847(p[792], s[878], c[864], s[879], c[879]);
fa fa848(p[823], s[879], c[865], s[880], c[880]);
fa fa849(p[854], s[880], c[866], s[881], c[881]);
fa fa850(p[885], s[881], c[867], s[882], c[882]);
fa fa851(p[916], s[882], c[868], s[883], c[883]);
fa fa852(p[947], s[883], c[869], s[884], c[884]);
fa fa853(p[978], s[884], c[870], s[885], c[885]);
fa fa854(p[1009], s[885], c[871], s[886], c[886]);

fa fa855(p[607], c[872], c[873], s[887], c[887]);
fa fa856(p[638], s[887], c[874], s[888], c[888]);
fa fa857(p[669], s[888], c[875], s[889], c[889]);
fa fa858(p[700], s[889], c[876], s[890], c[890]);
fa fa859(p[731], s[890], c[877], s[891], c[891]);
fa fa860(p[762], s[891], c[878], s[892], c[892]);
fa fa861(p[793], s[892], c[879], s[893], c[893]);
fa fa862(p[824], s[893], c[880], s[894], c[894]);
fa fa863(p[855], s[894], c[881], s[895], c[895]);
fa fa864(p[886], s[895], c[882], s[896], c[896]);
fa fa865(p[917], s[896], c[883], s[897], c[897]);
fa fa866(p[948], s[897], c[884], s[898], c[898]);
fa fa867(p[979], s[898], c[885], s[899], c[899]);
fa fa868(p[1010], s[899], c[886], s[900], c[900]);

fa fa869(p[639], c[887], c[888], s[901], c[901]);
fa fa870(p[670], s[901], c[889], s[902], c[902]);
fa fa871(p[701], s[902], c[890], s[903], c[903]);
fa fa872(p[732], s[903], c[891], s[904], c[904]);
fa fa873(p[763], s[904], c[892], s[905], c[905]);
fa fa874(p[794], s[905], c[893], s[906], c[906]);
fa fa875(p[825], s[906], c[894], s[907], c[907]);
fa fa876(p[856], s[907], c[895], s[908], c[908]);
fa fa877(p[887], s[908], c[896], s[909], c[909]);
fa fa878(p[918], s[909], c[897], s[910], c[910]);
fa fa879(p[949], s[910], c[898], s[911], c[911]);
fa fa880(p[980], s[911], c[899], s[912], c[912]);
fa fa881(p[1011], s[912], c[900], s[913], c[913]);

fa fa882(p[671], c[901], c[902], s[914], c[914]);
fa fa883(p[702], s[914], c[903], s[915], c[915]);
fa fa884(p[733], s[915], c[904], s[916], c[916]);
fa fa885(p[764], s[916], c[905], s[917], c[917]);
fa fa886(p[795], s[917], c[906], s[918], c[918]);
fa fa887(p[826], s[918], c[907], s[919], c[919]);
fa fa888(p[857], s[919], c[908], s[920], c[920]);
fa fa889(p[888], s[920], c[909], s[921], c[921]);
fa fa890(p[919], s[921], c[910], s[922], c[922]);
fa fa891(p[950], s[922], c[911], s[923], c[923]);
fa fa892(p[981], s[923], c[912], s[924], c[924]);
fa fa893(p[1012], s[924], c[913], s[925], c[925]);

fa fa894(p[703], c[914], c[915], s[926], c[926]);
fa fa895(p[734], s[926], c[916], s[927], c[927]);
fa fa896(p[765], s[927], c[917], s[928], c[928]);
fa fa897(p[796], s[928], c[918], s[929], c[929]);
fa fa898(p[827], s[929], c[919], s[930], c[930]);
fa fa899(p[858], s[930], c[920], s[931], c[931]);
fa fa900(p[889], s[931], c[921], s[932], c[932]);
fa fa901(p[920], s[932], c[922], s[933], c[933]);
fa fa902(p[951], s[933], c[923], s[934], c[934]);
fa fa903(p[982], s[934], c[924], s[935], c[935]);
fa fa904(p[1013], s[935], c[925], s[936], c[936]);

fa fa905(p[735], c[926], c[927], s[937], c[937]);
fa fa906(p[766], s[937], c[928], s[938], c[938]);
fa fa907(p[797], s[938], c[929], s[939], c[939]);
fa fa908(p[828], s[939], c[930], s[940], c[940]);
fa fa909(p[859], s[940], c[931], s[941], c[941]);
fa fa910(p[890], s[941], c[932], s[942], c[942]);
fa fa911(p[921], s[942], c[933], s[943], c[943]);
fa fa912(p[952], s[943], c[934], s[944], c[944]);
fa fa913(p[983], s[944], c[935], s[945], c[945]);
fa fa914(p[1014], s[945], c[936], s[946], c[946]);

fa fa915(p[767], c[937], c[938], s[947], c[947]);
fa fa916(p[798], s[947], c[939], s[948], c[948]);
fa fa917(p[829], s[948], c[940], s[949], c[949]);
fa fa918(p[860], s[949], c[941], s[950], c[950]);
fa fa919(p[891], s[950], c[942], s[951], c[951]);
fa fa920(p[922], s[951], c[943], s[952], c[952]);
fa fa921(p[953], s[952], c[944], s[953], c[953]);
fa fa922(p[984], s[953], c[945], s[954], c[954]);
fa fa923(p[1015], s[954], c[946], s[955], c[955]);

fa fa924(p[799], c[947], c[948], s[956], c[956]);
fa fa925(p[830], s[956], c[949], s[957], c[957]);
fa fa926(p[861], s[957], c[950], s[958], c[958]);
fa fa927(p[892], s[958], c[951], s[959], c[959]);
fa fa928(p[923], s[959], c[952], s[960], c[960]);
fa fa929(p[954], s[960], c[953], s[961], c[961]);
fa fa930(p[985], s[961], c[954], s[962], c[962]);
fa fa931(p[1016], s[962], c[955], s[963], c[963]);

fa fa932(p[831], c[956], c[957], s[964], c[964]);
fa fa933(p[862], s[964], c[958], s[965], c[965]);
fa fa934(p[893], s[965], c[959], s[966], c[966]);
fa fa935(p[924], s[966], c[960], s[967], c[967]);
fa fa936(p[955], s[967], c[961], s[968], c[968]);
fa fa937(p[986], s[968], c[962], s[969], c[969]);
fa fa938(p[1017], s[969], c[963], s[970], c[970]);

fa fa939(p[863], c[964], c[965], s[971], c[971]);
fa fa940(p[894], s[971], c[966], s[972], c[972]);
fa fa941(p[925], s[972], c[967], s[973], c[973]);
fa fa942(p[956], s[973], c[968], s[974], c[974]);
fa fa943(p[987], s[974], c[969], s[975], c[975]);
fa fa944(p[1018], s[975], c[970], s[976], c[976]);

fa fa945(p[895], c[971], c[972], s[977], c[977]);
fa fa946(p[926], s[977], c[973], s[978], c[978]);
fa fa947(p[957], s[978], c[974], s[979], c[979]);
fa fa948(p[988], s[979], c[975], s[980], c[980]);
fa fa949(p[1019], s[980], c[976], s[981], c[981]);

fa fa950(p[927], c[977], c[978], s[982], c[982]);
fa fa951(p[958], s[982], c[979], s[983], c[983]);
fa fa952(p[989], s[983], c[980], s[984], c[984]);
fa fa953(p[1020], s[984], c[981], s[985], c[985]);

fa fa954(p[959], c[982], c[983], s[986], c[986]);
fa fa955(p[990], s[986], c[984], s[987], c[987]);
fa fa956(p[1021], s[987], c[985], s[988], c[988]);

fa fa957(p[991], c[986], c[987], s[989], c[989]);
fa fa958(p[1022], s[989], c[988], s[990], c[990]);

fa fa959(p[1023], c[989], c[990], s[991], c[991]);

assign m[0] = p[0];
assign m[1] = s[0];
assign m[2] = s[2];
assign m[3] = s[5];
assign m[4] = s[9];
assign m[5] = s[14];
assign m[6] = s[20];
assign m[7] = s[27];
assign m[8] = s[35];
assign m[9] = s[44];
assign m[10] = s[54];
assign m[11] = s[65];
assign m[12] = s[77];
assign m[13] = s[90];
assign m[14] = s[104];
assign m[15] = s[119];
assign m[16] = s[135];
assign m[17] = s[152];
assign m[18] = s[170];
assign m[19] = s[189];
assign m[20] = s[209];
assign m[21] = s[230];
assign m[22] = s[252];
assign m[23] = s[275];
assign m[24] = s[299];
assign m[25] = s[324];
assign m[26] = s[350];
assign m[27] = s[377];
assign m[28] = s[405];
assign m[29] = s[434];
assign m[30] = s[464];
assign m[31] = s[495];
assign m[32] = s[526];
assign m[33] = s[556];
assign m[34] = s[585];
assign m[35] = s[613];
assign m[36] = s[640];
assign m[37] = s[666];
assign m[38] = s[691];
assign m[39] = s[715];
assign m[40] = s[738];
assign m[41] = s[760];
assign m[42] = s[781];
assign m[43] = s[801];
assign m[44] = s[820];
assign m[45] = s[838];
assign m[46] = s[855];
assign m[47] = s[871];
assign m[48] = s[886];
assign m[49] = s[900];
assign m[50] = s[913];
assign m[51] = s[925];
assign m[52] = s[936];
assign m[53] = s[946];
assign m[54] = s[955];
assign m[55] = s[963];
assign m[56] = s[970];
assign m[57] = s[976];
assign m[58] = s[981];
assign m[59] = s[985];
assign m[60] = s[988];
assign m[61] = s[990];
assign m[62] = s[991];
assign m[63] = c[991];

endmodule
