`timescale 1ns / 1ps
// Half Adder
module ha(input a, b,
    output sum, carry);
    assign sum = a ^ b;
    assign carry = a & b;
endmodule
// Full Adder
module fa (input a, b, cin,
    output sum, carry);
    assign sum = a ^ b ^ cin;
    assign carry =(a&b)|(b&cin)|(a&cin);
endmodule
module multi_16bit(
     input [15:0] A, B,
     output [31:0] P);
wire [255:0] p;
wire [239:0] s, c;
genvar i, j;// Generate Partial Products
  generate
    for(j = 0; j < 16; j = j + 1) begin: row
     for(i = 0; i < 16; i = i + 1) begin: col
      assign p[i + j*16] = A[i] & B[j];
     end
    end
  endgenerate
  
  

ha ha(p[1], p[16], s[0], c[0]);

fa fa0(p[2], p[17], c[0], s[1], c[1]);
ha ha1(p[32], s[1], s[2], c[2]);

fa fa1(p[3], p[18], c[1], s[3], c[3]);
fa fa2(p[33], s[3], c[2], s[4], c[4]);
ha ha2(p[48], s[4], s[5], c[5]);

fa fa3(p[4], p[19], c[3], s[6], c[6]);
fa fa4(p[34], s[6], c[4], s[7], c[7]);
fa fa5(p[49], s[7], c[5], s[8], c[8]);
ha ha3(p[64], s[8], s[9], c[9]);

fa fa6(p[5], p[120], c[6], s[10], c[10]);
fa fa7(p[35], s[10], c[7], s[11], c[11]);
fa fa8(p[50], s[11], c[8], s[12], c[12]);
fa fa9(p[65], s[12], c[9], s[13], c[13]);
ha ha4(p[80], s[13], s[14], c[14]);

fa fa10(p[6], p[21], c[10], s[15], c[15]);
fa fa11(p[36], s[15], c[11], s[16], c[16]);
fa fa12(p[51], s[16], c[12], s[17], c[17]);
fa fa13(p[66], s[17], c[13], s[18], c[18]);
fa fa14(p[81], s[18], c[14], s[19], c[19]);
ha ha5(p[96], s[19], s[20], c[20]);

fa fa15(p[7], p[22], c[15], s[21], c[21]);
fa fa16(p[37], s[21], c[16], s[22], c[22]);
fa fa17(p[52], s[22], c[17], s[23], c[23]);
fa fa18(p[67], s[23], c[18], s[24], c[24]);
fa fa19(p[82], s[24], c[19], s[25], c[25]);
fa fa20(p[97], s[25], c[20], s[26], c[26]);
ha ha6(p[112], s[26], s[27], c[27]);

fa fa21(p[8], p[23], c[21], s[28], c[28]);
fa fa22(p[38], s[28], c[22], s[29], c[29]);
fa fa23(p[53], s[29], c[23], s[30], c[30]);
fa fa24(p[68], s[30], c[24], s[31], c[31]);
fa fa25(p[83], s[31], c[25], s[32], c[32]);
fa fa26(p[98], s[32], c[26], s[33], c[33]);
fa fa27(p[113], s[33], c[27], s[34], c[34]);
ha ha7(p[128], s[34], s[35], c[35]);

fa fa28(p[9], p[24], c[28], s[36], c[36]);
fa fa29(p[39], s[36], c[29], s[37], c[37]);
fa fa30(p[54], s[37], c[30], s[38], c[38]);
fa fa31(p[69], s[38], c[31], s[39], c[39]);
fa fa32(p[84], s[39], c[32], s[40], c[40]);
fa fa33(p[99], s[40], c[33], s[41], c[41]);
fa fa34(p[114], s[41], c[34], s[42], c[42]);
fa fa35(p[129], s[42], c[35], s[43], c[43]);
ha ha8(p[144], s[43], s[44], c[44]);

fa fa36(p[10], p[25], c[36], s[45], c[45]);
fa fa37(p[40], s[45], c[37], s[46], c[46]);
fa fa38(p[55], s[46], c[38], s[47], c[47]);
fa fa39(p[70], s[47], c[39], s[48], c[48]);
fa fa40(p[85], s[48], c[40], s[49], c[49]);
fa fa41(p[100], s[49], c[41], s[50], c[50]);
fa fa42(p[115], s[50], c[42], s[51], c[51]);
fa fa43(p[130], s[51], c[43], s[52], c[52]);
fa fa44(p[145], s[52], c[44], s[53], c[53]);
ha ha9(p[160], s[53], s[54], c[54]);

fa fa45(p[11], p[26], c[45], s[55], c[55]);
fa fa46(p[41], s[55], c[46], s[56], c[56]);
fa fa47(p[56], s[56], c[47], s[57], c[57]);
fa fa48(p[71], s[57], c[48], s[58], c[58]);
fa fa49(p[86], s[58], c[49], s[59], c[59]);
fa fa50(p[101], s[59], c[50], s[60], c[60]);
fa fa51(p[116], s[60], c[51], s[61], c[61]);
fa fa52(p[131], s[61], c[52], s[62], c[62]);
fa fa53(p[146], s[62], c[53], s[63], c[63]);
fa fa54(p[161], s[63], c[54], s[64], c[64]);
ha ha10(p[176], s[64], s[65], c[65]);

fa fa55(p[12], p[27], c[55], s[66], c[66]);
fa fa56(p[42], s[66], c[56], s[67], c[67]);
fa fa57(p[57], s[67], c[57], s[68], c[68]);
fa fa58(p[72], s[68], c[58], s[69], c[69]);
fa fa59(p[87], s[69], c[59], s[70], c[70]);
fa fa60(p[102], s[70], c[60], s[71], c[71]);
fa fa61(p[117], s[71], c[61], s[72], c[72]);
fa fa62(p[132], s[72], c[62], s[73], c[73]);
fa fa63(p[147], s[73], c[63], s[74], c[74]);
fa fa64(p[162], s[74], c[64], s[75], c[75]);
fa fa65(p[177], s[75], c[65], s[76], c[76]);
ha ha11(p[192], s[76], s[77], c[77]);

fa fa66(p[13], p[28], c[66], s[78], c[78]);
fa fa67(p[43], s[78], c[67], s[79], c[79]);
fa fa68(p[58], s[79], c[68], s[80], c[80]);
fa fa69(p[73], s[80], c[69], s[81], c[81]);
fa fa70(p[88], s[81], c[70], s[82], c[82]);
fa fa71(p[103], s[82], c[71], s[83], c[83]);
fa fa72(p[118], s[83], c[72], s[84], c[84]);
fa fa73(p[133], s[84], c[73], s[85], c[85]);
fa fa74(p[148], s[85], c[74], s[86], c[86]);
fa fa75(p[163], s[86], c[75], s[87], c[87]);
fa fa76(p[178], s[87], c[76], s[88], c[88]);
fa fa77(p[193], s[88], c[77], s[89], c[89]);
ha ha12(p[208], s[89], s[90], c[90]);

fa fa78(p[14], p[29], c[78], s[91], c[91]);
fa fa79(p[44], s[91], c[79], s[92], c[92]);
fa fa80(p[59], s[92], c[80], s[93], c[93]);
fa fa81(p[74], s[93], c[81], s[94], c[94]);
fa fa82(p[89], s[94], c[82], s[95], c[95]);
fa fa83(p[104], s[95], c[83], s[96], c[96]);


fa fa84(p[119], s[96], c[84], s[97], c[97]);
fa fa85(p[134], s[97], c[85], s[98], c[98]);
fa fa86(p[149], s[98], c[86], s[99], c[99]);
fa fa87(p[164], s[99], c[87], s[100], c[100]);
fa fa88(p[179], s[100], c[88], s[101], c[101]);
fa fa89(p[194], s[101], c[89], s[102], c[102]);
fa fa90(p[209], s[102], c[90], s[103], c[103]);
ha ha13(p[224], s[103], s[104], c[104]);
fa fa91(p[15], p[30], c[91], s[105], c[105]);
fa fa92(p[45], s[105], c[92], s[106], c[106]);
fa fa93(p[60], s[106], c[93], s[107], c[107]);
fa fa94(p[75], s[107], c[94], s[108], c[108]);
fa fa95(p[90], s[108], c[95], s[109], c[109]);
fa fa96(p[105], s[109], c[96], s[110], c[110]);
fa fa97(p[120], s[110], c[97], s[111], c[111]);
fa fa98(p[135], s[111], c[98], s[112], c[112]);
fa fa99(p[150], s[112], c[99], s[113], c[113]);
fa fa100(p[165], s[113], c[100], s[114], c[114]);
fa fa101(p[180], s[114], c[101], s[115], c[115]);
fa fa102(p[195], s[115], c[102], s[116], c[116]);
fa fa103(p[210], s[116], c[103], s[117], c[117]);
fa fa104(p[225], s[117], c[104], s[118], c[118]);
ha ha14(p[240], s[118], s[119], c[119]);
fa fa105(p[31], c[105], c[106], s[120], c[120]);
fa fa106(p[46], s[120], c[107], s[121], c[121]);
fa fa107(p[61], s[121], c[108], s[122], c[122]);


fa fa108(p[76], s[122], c[109], s[123], c[123]);
fa fa109(p[91], s[123], c[110], s[124], c[124]);
fa fa110(p[106], s[124], c[111], s[125], c[125]);
fa fa111(p[121], s[125], c[112], s[126], c[126]);
fa fa112(p[136], s[126], c[113], s[127], c[127]);
fa fa113(p[151], s[127], c[114], s[128], c[128]);
fa fa114(p[166], s[128], c[115], s[129], c[129]);
fa fa115(p[181], s[129], c[116], s[130], c[130]);
fa fa116(p[196], s[130], c[117], s[131], c[131]);
fa fa117(p[211], s[131], c[118], s[132], c[132]);
fa fa118(p[226], s[132], c[119], s[133], c[133]);
ha ha15(p[241], s[133], s[134], c[134]);
fa fa119(p[47], c[120], c[121], s[135], c[135]);
fa fa121(p[62], s[135], c[122], s[136], c[136]);
fa fa122(p[77], s[136], c[123], s[137], c[137]);
fa fa123(p[92], s[137], c[124], s[138], c[138]);
fa fa124(p[107], s[138], c[125], s[139], c[139]);
fa fa125(p[122], s[139], c[126], s[140], c[140]);
fa fa126(p[137], s[140], c[127], s[141], c[141]);
fa fa127(p[152], s[141], c[128], s[142], c[142]);
fa fa128(p[167], s[142], c[129], s[143], c[143]);
fa fa129(p[182], s[143], c[130], s[144], c[144]);
fa fa130(p[197], s[144], c[131], s[145], c[145]);
fa fa131(p[212], s[145], c[132], s[146], c[146]);
fa fa132(p[227], s[146], c[133], s[147], c[147]);
fa fa133(p[242], s[147], c[134], s[148], c[148]);

fa fa134(p[63], c[135], c[136], s[149], c[149]);
fa fa135(p[78], s[149], c[137], s[150], c[150]);
fa fa136(p[93], s[150], c[138], s[151], c[151]);
fa fa137(p[108], s[151], c[139], s[152], c[152]);
fa fa138(p[123], s[152], c[140], s[153], c[153]);
fa fa139(p[138], s[153], c[141], s[154], c[154]);
fa fa140(p[153], s[154], c[142], s[155], c[155]);
fa fa141(p[168], s[155], c[143], s[156], c[156]);
fa fa142(p[183], s[156], c[144], s[157], c[157]);
fa fa143(p[198], s[157], c[145], s[158], c[158]);
fa fa144(p[213], s[158], c[146], s[159], c[159]);
fa fa145(p[228], s[159], c[147], s[160], c[160]);
fa fa146(p[243], s[160], c[148], s[161], c[161]);
fa fa147(p[79], c[149], c[150], s[162], c[162]);
fa fa148(p[94], s[162], c[151], s[163], c[163]);
fa fa149(p[109], s[163], c[152], s[164], c[164]);
fa fa150(p[124], s[164], c[153], s[165], c[165]);
fa fa151(p[139], s[165], c[154], s[166], c[166]);
fa fa152(p[154], s[166], c[155], s[167], c[167]);
fa fa153(p[169], s[167], c[156], s[168], c[168]);
fa fa154(p[184], s[168], c[157], s[169], c[169]);
fa fa155(p[199], s[169], c[158], s[170], c[170]);
fa fa156(p[214], s[170], c[159], s[171], c[171]);
fa fa157(p[229], s[171], c[160], s[172], c[172]);
fa fa158(p[244], s[172], c[161], s[173], c[173]);
fa fa159(p[95], c[162], c[163], s[174], c[174]);


fa fa160(p[110], s[174], c[164], s[175], c[175]);
fa fa161(p[125], s[175], c[165], s[176], c[176]);
fa fa162(p[140], s[176], c[166], s[177], c[177]);
fa fa163(p[155], s[177], c[167], s[178], c[178]);
fa fa164(p[170], s[178], c[168], s[179], c[179]);
fa fa165(p[185], s[179], c[169], s[180], c[180]);
fa fa166(p[200], s[180], c[170], s[181], c[181]);
fa fa167(p[215], s[181], c[171], s[182], c[182]);
fa fa168(p[230], s[182], c[172], s[183], c[183]);
fa fa169(p[245], s[183], c[173], s[184], c[184]);
fa fa170(p[111], c[174], c[175], s[185], c[185]);
fa fa171(p[126], s[185], c[176], s[186], c[186]);
fa fa172(p[141], s[186], c[177], s[187], c[187]);
fa fa173(p[156], s[187], c[178], s[188], c[188]);
fa fa174(p[171], s[188], c[179], s[189], c[189]);
fa fa175(p[186], s[189], c[180], s[190], c[190]);
fa fa176(p[201], s[190], c[181], s[191], c[191]);
fa fa177(p[216], s[191], c[182], s[192], c[192]);
fa fa178(p[231], s[192], c[183], s[193], c[193]);
fa fa179(p[246], s[193], c[184], s[194], c[194]);
fa fa180(p[127], c[185], c[186], s[195], c[195]);
fa fa181(p[142], s[195], c[187], s[196], c[196]);
fa fa182(p[157], s[196], c[188], s[197], c[197]);
fa fa183(p[172], s[197], c[189], s[198], c[198]);
fa fa184(p[187], s[198], c[190], s[199], c[199]);
fa fa185(p[202], s[199], c[191], s[200], c[200]);

fa fa186(p[217], s[200], c[192], s[201], c[201]);
fa fa187(p[232], s[201], c[193], s[202], c[202]);
fa fa188(p[247], s[202], c[194], s[203], c[203]);
fa fa189(p[143], c[195], c[196], s[204], c[204]);
fa fa190(p[158], s[204], c[197], s[205], c[205]);
fa fa191(p[173], s[205], c[198], s[206], c[206]);
fa fa192(p[188], s[206], c[199], s[207], c[207]);
fa fa193(p[203], s[207], c[200], s[208], c[208]);
fa fa194(p[218], s[208], c[201], s[209], c[209]);
fa fa195(p[233], s[209], c[202], s[210], c[210]);
fa fa196(p[248], s[210], c[203], s[211], c[211]);
fa fa197(p[159], c[204], c[205], s[212], c[212]);
fa fa198(p[174], s[212], c[206], s[213], c[213]);
fa fa199(p[189], s[213], c[207], s[214], c[214]);
fa fa200(p[204], s[214], c[208], s[215], c[215]);
fa fa201(p[219], s[215], c[209], s[216], c[216]);
fa fa202(p[234], s[216], c[210], s[217], c[217]);
fa fa203(p[249], s[217], c[211], s[218], c[218]);
fa fa204(p[175], c[212], c[213], s[219], c[219]);
fa fa205(p[190], s[219], c[214], s[220], c[220]);
fa fa206(p[205], s[220], c[215], s[221], c[221]);
fa fa207(p[220], s[221], c[216], s[222], c[222]);
fa fa208(p[235], s[222], c[217], s[223], c[223]);
fa fa209(p[250], s[223], c[218], s[224], c[224]);
fa fa210(p[191], c[219], c[220], s[225], c[225]);
fa fa211(p[206], s[225], c[221], s[226], c[226]);

fa fa212(p[221], s[226], c[222], s[227], c[227]);
fa fa213(p[236], s[227], c[223], s[228], c[228]);
fa fa214(p[251], s[228], c[224], s[229], c[229]);
fa fa215(p[207], c[225], c[226], s[230], c[230]);
fa fa216(p[222], s[230], c[227], s[231], c[231]);
fa fa217(p[237], s[231], c[228], s[232], c[232]);
fa fa218(p[252], s[232], c[229], s[233], c[233]);
fa fa219(p[223], c[230], c[231], s[234], c[234]);
fa fa220(p[238], s[234], c[232], s[235], c[235]);
fa fa221(p[253], s[235], c[233], s[236], c[236]);
fa fa222(p[239], c[234], c[235], s[237], c[237]);
fa fa223(p[254], s[237], c[236], s[238], c[238]);
fa fa224(p[255], c[237], c[238], s[239], c[239]);
assign P[0] = p[0];
assign P[1] = s[0];
assign P[2] = s[2];
assign P[3] = s[5];
assign P[4] = s[9];
assign P[5] = s[14];
assign P[6] = s[20];
assign P[7] = s[27];
assign P[8] = s[35];
assign P[9] = s[44];
assign P[10] = s[54];


assign P[11] = s[65];
assign P[12] = s[77];
assign P[13] = s[90];
assign P[14] = s[104];
assign P[15] = s[119];
assign P[16] = s[134];
assign P[17] = s[148];
assign P[18] = s[161];
assign P[19] = s[173];
assign P[20] = s[184];
assign P[21] = s[194];
assign P[22] = s[203];
assign P[23] = s[211];
assign P[24] = s[218];
assign P[25] = s[224];
assign P[26] = s[229];
assign P[27] = s[233];
assign P[28] = s[236];
assign P[29] = s[238];
assign P[30] = s[239];
assign P[31] = c[239];
endmodule
